library ieee;
use ieee.std_logic_1164.all;

entity four_second_timer is
	port (
		a: in std_ulogic;
		b: out std_ulogic;
	);
	
end entity four_second_timer;

architecture count of four_second_timer is

begin
	
end architecture count;
